//-- EE 2019

module	greenwinBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
);
// generating a green wining screen bitmap 

localparam  int OBJECT_HEIGHT_Y = 64;
localparam  int OBJECT_WIDTH_X = 64;

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 


logic [0:OBJECT_WIDTH_X-1] [0:OBJECT_HEIGHT_Y-1] [8-1:0] object_colors = {
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h35, 8'h35, 8'h15, 8'h35, 8'h35, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h35, 8'h15, 8'h35, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'hBA, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h5A, 8'hFF, 8'hFF, 8'h55, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'h55, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h15, 8'h35, 8'hBA, 8'hBA, 8'hBA, 8'h35, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hBA, 8'hBA, 8'h7A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h5A, 8'h15, 8'h35, 8'h9A, 8'hBA, 8'hBA, 8'hBA, 8'hBA, 8'hBA, 8'hFF, 8'hFF, 8'hDF, 8'h35, 8'h15, 8'h5A, 8'hBA, 8'hBA, 8'hBA, 8'hBA, 8'hBA, 8'hDF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h35, 8'h35, 8'h9A, 8'hFF, 8'h5A, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'h11F, 8'h11F, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h5A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h15, 8'h55, 8'hFF, 8'h55, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h5A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h15, 8'h15, 8'hDF, 8'h56, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hDF, 8'hDF, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h5A, 8'h15, 8'h35, 8'hBA, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h35, 8'h15, 8'h5A, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h35, 8'h35, 8'h15, 8'h9A, 8'h7A, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h15, 8'h35, 8'hFF, 8'h9A, 8'h15, 8'h35, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'hBA, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h35, 8'h15, 8'h55, 8'h56, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h55, 8'hFF, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h15, 8'h35, 8'hFF, 8'h9A, 8'h15, 8'h35, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'hBA, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h7A, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h35, 8'hDF, 8'hDF, 8'hBA, 8'h35, 8'h35, 8'h55, 8'hFF, 8'hFF, 8'hBA, 8'h35, 8'h35, 8'h7A, 8'hBF, 8'hBF, 8'h9A, 8'h35, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h5A, 8'h15, 8'h35, 8'hBA, 8'hBB, 8'hBB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h35, 8'h35, 8'h5A, 8'hBF, 8'hBA, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h35, 8'hBA, 8'h35, 8'h35, 8'h35, 8'h35, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h5A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'hDF, 8'h5A, 8'h15, 8'h35, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h5A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'hDF, 8'hBA, 8'h15, 8'h15, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h35, 8'hBA, 8'hDF, 8'hBF, 8'h35, 8'h15, 8'h55, 8'hFF, 8'hFF, 8'hBA, 8'h35, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h5A, 8'h15, 8'h35, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'h35, 8'h15, 8'h5A, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'h35, 8'h35, 8'h35, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h15, 8'h35, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'hBF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'hBF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'hBF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hBF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBF, 8'hBF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hBF, 8'hBF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hBF, 8'hDF, 8'hDF, 8'hBF, 8'hDF, 8'hDF, 8'hBF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hBF, 8'hBF, 8'hDF, 8'hDF, 8'hBF, 8'hDF, 8'hDF, 8'hBF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hBF, 8'hBF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hBF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h5A, 8'h5A, 8'h9A, 8'hFF, 8'hFF, 8'hBB, 8'h5A, 8'h5A, 8'hBA, 8'hFF, 8'hFF, 8'hBA, 8'h5A, 8'h5A, 8'hBB, 8'hFF, 8'hFF, 8'h7A, 8'h5A, 8'h7A, 8'h7A, 8'h5A, 8'h7A, 8'h7A, 8'h5A, 8'h7A, 8'hFF, 8'hFF, 8'hDF, 8'h5A, 8'h5A, 8'h9A, 8'hFF, 8'hFF, 8'hBB, 8'h5A, 8'h5A, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h00, 8'h55, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'hFF, 8'h7A, 8'hFF, 8'hFF, 8'h7A, 8'h00, 8'h15, 8'hBB, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'h9A, 8'hFF, 8'hFF, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h55, 8'hFF, 8'hFF, 8'h55, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h15, 8'hBA, 8'h11F, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'h56, 8'h15, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'h55, 8'h15, 8'h55, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h55, 8'h5A, 8'h35, 8'h15, 8'h35, 8'h5A, 8'h56, 8'h7A, 8'hFF, 8'hFF, 8'hBB, 8'h15, 8'h15, 8'h35, 8'h7A, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'hBA, 8'hDF, 8'h35, 8'h15, 8'h15, 8'h35, 8'hBF, 8'hDF, 8'h35, 8'h15, 8'h5A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h35, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'h15, 8'h9A, 8'hDF, 8'h35, 8'h15, 8'h15, 8'h15, 8'h9A, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h15, 8'hBA, 8'hBA, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h7A, 8'hBA, 8'h35, 8'h15, 8'h15, 8'h35, 8'h7A, 8'h9A, 8'h35, 8'h15, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h15, 8'h5A, 8'hBA, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h35, 8'h35, 8'h56, 8'h7A, 8'h35, 8'h35, 8'h35, 8'h35, 8'h7A, 8'h7A, 8'h35, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBB, 8'h35, 8'h35, 8'h35, 8'h35, 8'h35, 8'h9A, 8'h35, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'h35, 8'h15, 8'h15, 8'h15, 8'h35, 8'h35, 8'h35, 8'h15, 8'h15, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h55, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5A, 8'h15, 8'h15, 8'h15, 8'h35, 8'h35, 8'h35, 8'h35, 8'h15, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h55, 8'h15, 8'h15, 8'h35, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'h35, 8'h35, 8'h35, 8'h35, 8'h5A, 8'h7A, 8'h35, 8'h35, 8'h35, 8'h35, 8'h7A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBB, 8'h35, 8'h15, 8'h7A, 8'h5A, 8'h35, 8'h35, 8'h35, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h15, 8'h35, 8'h7A, 8'h9A, 8'h35, 8'h15, 8'h15, 8'h35, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'h9A, 8'h15, 8'h35, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h15, 8'h15, 8'h15, 8'h15, 8'h9A, 8'hBA, 8'h15, 8'h15, 8'h15, 8'h15, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hDF, 8'h15, 8'h35, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h35, 8'h15, 8'h15, 8'h35, 8'hBB, 8'hDF, 8'h35, 8'h15, 8'h15, 8'h35, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'h56, 8'h35, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5A, 8'h35, 8'h35, 8'h35, 8'hDF, 8'hFF, 8'h56, 8'h35, 8'h35, 8'h55, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h55, 8'h56, 8'h35, 8'h35, 8'h35, 8'h56, 8'h55, 8'h7A, 8'hFF, 8'hFF, 8'hBB, 8'h35, 8'h15, 8'h7A, 8'h11F, 8'h9A, 8'h35, 8'h35, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'h5A, 8'h15, 8'h15, 8'h56, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'h15, 8'h7A, 8'hFF, 8'hDF, 8'h35, 8'h15, 8'h15, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'h15, 8'hFF, 8'h5A, 8'hFF, 8'hFF, 8'h7A, 8'hFF, 8'hFF, 8'h7A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h35, 8'hFF, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h35, 8'hFF, 8'hFF, 8'hBA, 8'h15, 8'hFF, 8'h7A, 8'hFF, 8'hFF, 8'h5A, 8'h15, 8'hFF, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h7A, 8'h5A, 8'hBA, 8'hFF, 8'hFF, 8'hBA, 8'h5A, 8'h5A, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'h5A, 8'h7A, 8'h7A, 8'h7A, 8'h7A, 8'h7A, 8'h7A, 8'h7A, 8'hFF, 8'hFF, 8'hDF, 8'h7A, 8'h5A, 8'h9A, 8'hFF, 8'hFF, 8'hBA, 8'h5A, 8'h5A, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF }
};


// pipeline (ff) to get the pixel color from the array 	 

//======--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		if (InsideRectangle == 1'b1 )  // inside an external bracket 
			RGBout <= object_colors[offsetY/4][offsetX/4];	//get RGB from the colors table  
		else 
			RGBout <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
	end 
end

//======--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   

endmodule