

module strong_matrix_init	(	//this module creat 4 difrent maps of bricks and send them to the square
					output	logic	[0:14] [0:19]		mat_out0,
					output	logic	[0:14] [0:19]		mat_out1,
					output	logic	[0:14] [0:19]		mat_out2,
					output	logic	[0:14] [0:19]		mat_out3
);

//15 lines of y
//20 lines of x

bit [0:14] [0:19] mat0  = 


{
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,

};
bit [0:14] [0:19] mat1  = 


{
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h1,	1'h1,	1'h1,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h1,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h1,	1'h1,	1'h1,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h1,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h1,	1'h1,	1'h1,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h1,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h1,	1'h1,	1'h1,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h1,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,


};
bit [0:14] [0:19] mat2  = 


{
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,


};
bit [0:14] [0:19] mat3  = 


{
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h1,	1'h1,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,	1'h0,
};															
 
																	
	assign mat_out0 = mat0 ;
	assign mat_out1 = mat1 ;
	assign mat_out2 = mat2 ;
	assign mat_out3 = mat3 ;

endmodule